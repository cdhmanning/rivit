/*
 *
 */

typedef logic [xreg_width - 1 : 0] xreg_t;
